module alu(input [31:0] A,
           input [31:0] B, 
           input [ 2:0] ALUOp,
           output Z, // Z = 1, if Result = 0
           output V, // V = 1, if Overflow
           output C //  C32 = 1, if Carry-Out
           output [31:0] Result);

           




endmodule